module mycpu_top(
    input  aclk   ,
    input  aresetn,
    // read req channel
    output [ 3:0] arid   , // 读请求ID
    output [31:0] araddr , // 读请求地址
    output [ 7:0] arlen  , // 读请求传输长度（数据传输拍数）
    output [ 2:0] arsize , // 读请求传输大小（数据传输每拍的字节数）
    output [ 1:0] arburst, // 传输类型
    output [ 1:0] arlock , // 原子锁
    output [ 3:0] arcache, // Cache属性
    output [ 2:0] arprot , // 保护属性
    output        arvalid, // 读请求地址有效
    input         arready, // 读请求地址握手信号
    // read response channel
    input [ 3:0]  rid    , // 读请求ID号，同一请求rid与arid一致
    input [31:0]  rdata  , // 读请求读出的数据
    input [ 1:0]  rresp  , // 读请求是否完成
    input         rlast  , // 读请求最后一拍数据的指示信号
    input         rvalid , // 读请求数据有效
    output        rready , // Master端准备好接受数据
    // write req channel
    output [ 3:0] awid   , // 写请求的ID号
    output [31:0] awaddr , // 写请求的地址
    output [ 7:0] awlen  , // 写请求传输长度（拍数）
    output [ 2:0] awsize , // 写请求传输每拍字节数
    output [ 1:0] awburst, // 写请求传输类型
    output [ 1:0] awlock , // 原子锁
    output [ 3:0] awcache, // Cache属性
    output [ 2:0] awprot , // 保护属性
    output        awvalid, // 写请求地址有效
    input         awready, // Slave端准备好接受地址传输   
    // write data channel
    output [ 3:0] wid    , // 写请求的ID号
    output [31:0] wdata  , // 写请求的写数据
    output [ 3:0] wstrb  , // 写请求字节选通位
    output        wlast  , // 写请求的最后一拍数据的指示信号
    output        wvalid , // 写数据有效
    input         wready , // Slave端准备好接受写数据传输   
    // write response channel
    input  [ 3:0] bid    , // 写请求的ID号
    input  [ 1:0] bresp  , // 写请求完成信号
    input         bvalid , // 写请求响应有效
    output        bready , // Master端准备好接收响应信号
    // trace debug interface
    output wire [31:0] debug_wb_pc,
    output wire [ 3:0] debug_wb_rf_we,
    output wire [ 4:0] debug_wb_rf_wnum,
    output wire [31:0] debug_wb_rf_wdata
);

    // inst sram interface (some signals modified due to I-Cache)
    wire        inst_sram_req;
    wire        inst_sram_wr;
    wire [ 1:0] inst_sram_size;
    wire [ 3:0] inst_sram_wstrb;
    wire [31:0] inst_sram_addr;
    wire [31:0] inst_sram_wdata;
    wire        icache_cpu_addr_ok;
    wire        icache_cpu_data_ok;
    wire [31:0] icache_cpu_rdata;
    // data sram interface
    wire        data_sram_req;
    wire        data_sram_wr;
    wire [ 1:0] data_sram_size;
    wire [ 3:0] data_sram_wstrb;
    wire [31:0] data_sram_addr;
    wire [31:0] data_sram_wdata;
    wire        data_sram_addr_ok;
    wire        data_sram_data_ok;
    wire [31:0] data_sram_rdata;
    // I-Cache interface 
    wire         icache_axi_rd_req;
    wire [  2:0] icache_axi_rd_type;
    wire [ 31:0] icache_axi_rd_addr;
    wire         icache_axi_rd_rdy;
	wire         icache_axi_ret_valid;
	wire         icache_axi_ret_last;
	wire [ 31:0] icache_axi_ret_data;
    // wr_* signals reserved to avoid ports suspending
    wire         icache_axi_wr_req;
    wire [  2:0] icache_axi_wr_type;
    wire [ 31:0] icache_axi_wr_addr;
	wire [  3:0] icache_axi_wr_wstrb;
    wire [127:0] icache_wr_data;

    mycpu_core my_core(
        .clk            (aclk       ),
        .resetn         (aresetn    ),
        // inst sram interface
        .inst_sram_req      (inst_sram_req      ),
        .inst_sram_wr       (inst_sram_wr       ),
        .inst_sram_size     (inst_sram_size     ),
        .inst_sram_wstrb    (inst_sram_wstrb    ),
        .inst_sram_addr     (inst_sram_addr     ),
        .inst_sram_wdata    (inst_sram_wdata    ),
        .inst_sram_addr_ok  (icache_cpu_addr_ok ),
        .inst_sram_data_ok  (icache_cpu_data_ok ),
        .inst_sram_rdata    (icache_cpu_rdata   ),
        // data sram interface
        .data_sram_req      (data_sram_req      ),
        .data_sram_wr       (data_sram_wr       ),
        .data_sram_size     (data_sram_size     ),
        .data_sram_wstrb    (data_sram_wstrb    ),
        .data_sram_addr     (data_sram_addr     ),
        .data_sram_wdata    (data_sram_wdata    ),
        .data_sram_addr_ok  (data_sram_addr_ok  ),
        .data_sram_data_ok  (data_sram_data_ok  ),
        .data_sram_rdata    (data_sram_rdata    ),
        // trace debug interface
        .debug_wb_pc        (debug_wb_pc        ),
        .debug_wb_rf_we     (debug_wb_rf_we     ),
        .debug_wb_rf_wnum   (debug_wb_rf_wnum   ),
        .debug_wb_rf_wdata  (debug_wb_rf_wdata  )
    );

    cache my_icache(
        .clk      (aclk                 ),
        .resetn   (aresetn              ),
        // cpu-icache interface
        .valid    (inst_sram_req        ),
	    .op       (inst_sram_wr         ),
        .index    (inst_sram_addr[11:4] ),
	    .tag      (inst_sram_addr[31:12]),
	    .offset   (inst_sram_addr[3:0]  ),
        .wstrb    (inst_sram_wstrb      ),
	    .wdata    (inst_sram_wdata      ),
	    .addr_ok  (icache_cpu_addr_ok   ),
	    .data_ok  (icache_cpu_data_ok   ),
	    .rdata    (icache_cpu_rdata     ),
	    // icache-axi interface
        .rd_req   (icache_axi_rd_req    ),
        .rd_type  (icache_axi_rd_type   ),
        .rd_addr  (icache_axi_rd_addr   ),
	    .rd_rdy   (icache_axi_rd_rdy    ),
	    .ret_valid(icache_axi_ret_valid ),
	    .ret_last (icache_axi_ret_last  ),
	    .ret_data (icache_axi_ret_data  ),
        // invalid in I-Cache (reserved to avoid ports suspending)
        .wr_req   (icache_axi_wr_req    ),
        .wr_type  (icache_axi_wr_type   ),
        .wr_addr  (icache_axi_wr_addr   ),
	    .wr_wstrb (icache_axi_wr_wstrb  ),
        .wr_data  (icache_wr_data       ),
	    .wr_rdy   (1'b1                 )
    );

    bridge_sram_axi my_bridge_sram_axi(
        .aclk               (aclk               ),
        .aresetn            (aresetn            ),

        .arid               (arid               ),
        .araddr             (araddr             ),
        .arlen              (arlen              ),
        .arsize             (arsize             ),
        .arburst            (arburst            ),
        .arlock             (arlock             ),
        .arcache            (arcache            ),
        .arprot             (arprot             ),
        .arvalid            (arvalid            ),
        .arready            (arready            ),

        .rid                (rid                ),
        .rdata              (rdata              ),
        .rvalid             (rvalid             ),
        .rlast              (rlast              ),
        .rready             (rready             ),
        .rresp              (rresp              ),

        .awid               (awid               ),
        .awaddr             (awaddr             ),
        .awlen              (awlen              ),
        .awsize             (awsize             ),
        .awburst            (awburst            ),
        .awlock             (awlock             ),
        .awcache            (awcache            ),
        .awprot             (awprot             ),
        .awvalid            (awvalid            ),
        .awready            (awready            ),

        .wid                (wid                ),
        .wdata              (wdata              ),
        .wstrb              (wstrb              ),
        .wlast              (wlast              ),
        .wvalid             (wvalid             ),
        .wready             (wready             ),

        .bid                (bid                ),
        .bvalid             (bvalid             ),
        .bready             (bready             ),
        .bresp              (bresp              ),
        // modified due to I-Cache
        .icache_axi_rd_req   (icache_axi_rd_req   ),
        .icache_axi_rd_type  (icache_axi_rd_type  ),
        .icache_axi_rd_addr  (icache_axi_rd_addr  ),
	    .icache_axi_rd_rdy   (icache_axi_rd_rdy   ),
	    .icache_axi_ret_valid(icache_axi_ret_valid),
	    .icache_axi_ret_last (icache_axi_ret_last ),
	    .icache_axi_ret_data (icache_axi_ret_data ),

        .data_sram_req      (data_sram_req      ),
        .data_sram_wr       (data_sram_wr       ),
        .data_sram_size     (data_sram_size     ),
        .data_sram_addr     (data_sram_addr     ),
        .data_sram_wstrb    (data_sram_wstrb    ),
        .data_sram_wdata    (data_sram_wdata    ),
        .data_sram_addr_ok  (data_sram_addr_ok  ),
        .data_sram_data_ok  (data_sram_data_ok  ),
        .data_sram_rdata    (data_sram_rdata    )
    );

endmodule
